import uvm_pkg::*;
`include "uvm_macros.svh"

class fc_env extends uvm_env;
endclass: fc_env