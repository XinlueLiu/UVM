`define NUM_CNT_BITS 4